library verilog;
use verilog.vl_types.all;
entity wrong_code_tester_vlg_vec_tst is
end wrong_code_tester_vlg_vec_tst;
