LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY Mux IS
	PORT (
		-- Input ports
		A1 : IN STD_LOGIC_VECTOR(6 downto 0);
		A2 : IN STD_LOGIC_VECTOR(6 downto 0);
		A3 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		A4 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		B1 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		B2 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		B3 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		B4 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		B5 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		B6 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		VIEW   : IN std_LOGIC;
		-- Output ports
		C1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		C2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		C3 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		C4 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		C5 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		C6 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END Mux;

ARCHITECTURE Mux_impl OF Mux IS
BEGIN

	PROCESS (A1,A2,A3,A4,B1,B2,B3,B4,B5,B6) IS
		-- Declaration(s) 
	BEGIN
		IF VIEW = '0' THEN
			
			C1 <= "1111111";
			C2 <= "1111111";
			C3 <= A1;
			C4 <= A2;
			C5 <= A3;
			C6 <= A4;
		else
			C1 <= B1;
			C2 <= B2;
			C3 <= B3;
			C4 <= B4;
			C5 <= B5;
			C6 <= B6;

		END IF;
	END PROCESS;
END Mux_impl;