library verilog;
use verilog.vl_types.all;
entity Code_lock_vlg_vec_tst is
end Code_lock_vlg_vec_tst;
