--LIBRARY ieee;
--USE ieee.std_logic_1164.ALL;
--USE ieee.numeric_std.ALL;
--USE work.ALL;
--
--ENTITY demux_tester IS
--	PORT
--	(
--		-- Input ports
--		SW     : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
--		KEY    : in STD_LOGIC_VECTOR(1 DOWNTO 0);
--
--		-- Output ports
--		HEX0   : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
--		HEX1   : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
--		HEX2   : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
--
--	);
--END demux_tester;
--
--ARCHITECTURE demux_tester_impl OF demux_tester IS
--BEGIN
--
--	
--
--
--END demux_tester_impl;